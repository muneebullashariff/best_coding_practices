Always use the branch to do the development work and once everything works on the development-branch go ahead and merge the changes
into the master-branch. DON'T MESS WITH THE MASTER

Please refer the article below as how to achieve this:
https://thenewstack.io/dont-mess-with-the-master-working-with-branches-in-git-and-github/
