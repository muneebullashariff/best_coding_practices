`ifndef _<<USER_FILENAME>>_INCLUDED_
`define _<<USER_FILENAME>>_INCLUDED_

//--------------------------------------------------------------------------------------------
// Class: <<user_classname>> 
// <Description_here>
//--------------------------------------------------------------------------------------------
class <<user_classname>> extends uvm_component;
  `uvm_component_utils(<<user_classname>>)

  //-------------------------------------------------------
  //Externally defined Tasks and Functions 
  //-------------------------------------------------------
  extern function new(string name = "<<user_classname>>", uvm_component parent = null);
  extern virtual function void build_phase(uvm_phase phase);
  extern virtual function void connect_phase(uvm_phase phase);
  extern virtual function void end_of_elaboration_phase(uvm_phase phase);
  extern virtual function void start_of_simulation_phase(uvm_phase phase);
  extern virtual task run_phase(uvm_phase phase);

endclass: <<user_classname>>

//--------------------------------------------------------------------------------------------
// Construct: new
// 
// Parameters:
//  name - <<user_classname>>
//  parent - parent under which this component is created
//--------------------------------------------------------------------------------------------
function <<user_classname>>::new(string name = "<<user_classname>>",      
                                 uvm_component parent = null);
  super.new(name, parent);
endfunction: new

//--------------------------------------------------------------------------------------------
// Function: build_phase
// <Description_here>
//
// Parameters:
//  phase - uvm phase
//--------------------------------------------------------------------------------------------
function void <<user_classname>>::build_phase(uvm_phase phase);
  super.build_phase(phase);
endfunction: build_phase

//--------------------------------------------------------------------------------------------
// Function: connect_phase
// <Description_here>
//
// Parameters:
//  phase - uvm phase
//--------------------------------------------------------------------------------------------
function void <<user_classname>>::connect_phase(uvm_phase phase);
  super.connect_phase(phase);
endfunction: connect_phase

//--------------------------------------------------------------------------------------------
// Function: end_of_elaboration_phase
// <Description_here>
//
// Parameters:
//  phase - uvm phase
//--------------------------------------------------------------------------------------------
function void <<user_classname>>::end_of_elaboration_phase(uvm_phase phase);
  super.end_of_elaboration_phase(phase);
endfunction: end_of_elaboration_phase

//--------------------------------------------------------------------------------------------
// Function: start_of_simulation_phase
// <Description_here>
//
// Parameters:
//  phase - uvm phase
//--------------------------------------------------------------------------------------------
function void <<user_classname>>::start_of_simulation_phase(uvm_phase phase);
  super.start_of_simulation_phase(phase);
endfunction: start_of_simulation_phase

//--------------------------------------------------------------------------------------------
// Task: run_phase
// <Description_here>
// 
// Parameters: 
//  phase - uvm phase
//--------------------------------------------------------------------------------------------
task <<user_classname>>::run_phase(uvm_phase phaase);

  phase.raise_objection(this, "<<user_classname>>");

  super.run_phase(phase);

  // Work here
  // ...

  phase.drop_objection(this);

endtask: run_phase

`endif
